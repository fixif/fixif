--*********testbench*********--
---testbench---

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use work.all;

entity test is 
end;

architecture tb of test is
  component top_cell
    port(
     i0 : IN std_logic_vector (15 downto 0);
     i1 : IN std_logic_vector (15 downto 0);
     i2 : IN std_logic_vector (15 downto 0);
     i3 : IN std_logic_vector (15 downto 0);
     oo : OUT std_logic_vector (15 downto 0)
  );
  end component;
  signal i0 : std_logic_vector (15 downto 0) := x"0000";
  signal i1 : std_logic_vector (15 downto 0) := x"0000";
  signal i2 : std_logic_vector (15 downto 0) := x"0000";
  signal i3 : std_logic_vector (15 downto 0) := x"0000";
  signal oo : std_logic_vector(15 downto 0);

  begin
    instance : entity work.top_cell port map(i0 => i0,i1 => i1,i2 => i2,i3 => i3,oo => oo);

    simu : process is
    begin
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0000";
      i2<=x"0000";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0000";
      i2<=x"0000";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0000";
      i2<=x"0000";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0000";
      i2<=x"0000";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0000";
      i2<=x"0001";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0000";
      i2<=x"0001";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0000";
      i2<=x"0001";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0000";
      i2<=x"0001";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0000";
      i2<=x"0002";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0000";
      i2<=x"0002";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0000";
      i2<=x"0002";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0000";
      i2<=x"0002";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0000";
      i2<=x"0003";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0000";
      i2<=x"0003";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0000";
      i2<=x"0003";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0000";
      i2<=x"0003";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0001";
      i2<=x"0000";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0001";
      i2<=x"0000";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0001";
      i2<=x"0000";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0001";
      i2<=x"0000";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0001";
      i2<=x"0001";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0001";
      i2<=x"0001";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0001";
      i2<=x"0001";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0001";
      i2<=x"0001";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0001";
      i2<=x"0002";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0001";
      i2<=x"0002";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0001";
      i2<=x"0002";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0001";
      i2<=x"0002";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0001";
      i2<=x"0003";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0001";
      i2<=x"0003";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0001";
      i2<=x"0003";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0001";
      i2<=x"0003";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0002";
      i2<=x"0000";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0002";
      i2<=x"0000";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0002";
      i2<=x"0000";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0002";
      i2<=x"0000";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0002";
      i2<=x"0001";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0002";
      i2<=x"0001";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0002";
      i2<=x"0001";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0002";
      i2<=x"0001";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0002";
      i2<=x"0002";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0002";
      i2<=x"0002";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0002";
      i2<=x"0002";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0002";
      i2<=x"0002";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0002";
      i2<=x"0003";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0002";
      i2<=x"0003";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0002";
      i2<=x"0003";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0002";
      i2<=x"0003";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0003";
      i2<=x"0000";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0003";
      i2<=x"0000";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0003";
      i2<=x"0000";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0003";
      i2<=x"0000";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0003";
      i2<=x"0001";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0003";
      i2<=x"0001";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0003";
      i2<=x"0001";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0003";
      i2<=x"0001";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0003";
      i2<=x"0002";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0003";
      i2<=x"0002";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0003";
      i2<=x"0002";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0003";
      i2<=x"0002";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0003";
      i2<=x"0003";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0003";
      i2<=x"0003";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0003";
      i2<=x"0003";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0000";
      i1<=x"0003";
      i2<=x"0003";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0000";
      i2<=x"0000";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0000";
      i2<=x"0000";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0000";
      i2<=x"0000";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0000";
      i2<=x"0000";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0000";
      i2<=x"0001";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0000";
      i2<=x"0001";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0000";
      i2<=x"0001";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0000";
      i2<=x"0001";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0000";
      i2<=x"0002";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0000";
      i2<=x"0002";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0000";
      i2<=x"0002";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0000";
      i2<=x"0002";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0000";
      i2<=x"0003";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0000";
      i2<=x"0003";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0000";
      i2<=x"0003";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0000";
      i2<=x"0003";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0001";
      i2<=x"0000";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0001";
      i2<=x"0000";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0001";
      i2<=x"0000";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0001";
      i2<=x"0000";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0001";
      i2<=x"0001";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0001";
      i2<=x"0001";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0001";
      i2<=x"0001";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0001";
      i2<=x"0001";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0001";
      i2<=x"0002";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0001";
      i2<=x"0002";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0001";
      i2<=x"0002";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0001";
      i2<=x"0002";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0001";
      i2<=x"0003";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0001";
      i2<=x"0003";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0001";
      i2<=x"0003";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0001";
      i2<=x"0003";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0002";
      i2<=x"0000";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0002";
      i2<=x"0000";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0002";
      i2<=x"0000";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0002";
      i2<=x"0000";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0002";
      i2<=x"0001";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0002";
      i2<=x"0001";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0002";
      i2<=x"0001";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0002";
      i2<=x"0001";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0002";
      i2<=x"0002";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0002";
      i2<=x"0002";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0002";
      i2<=x"0002";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0002";
      i2<=x"0002";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0002";
      i2<=x"0003";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0002";
      i2<=x"0003";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0002";
      i2<=x"0003";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0002";
      i2<=x"0003";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0003";
      i2<=x"0000";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0003";
      i2<=x"0000";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0003";
      i2<=x"0000";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0003";
      i2<=x"0000";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0003";
      i2<=x"0001";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0003";
      i2<=x"0001";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0003";
      i2<=x"0001";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0003";
      i2<=x"0001";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0003";
      i2<=x"0002";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0003";
      i2<=x"0002";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0003";
      i2<=x"0002";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0003";
      i2<=x"0002";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0003";
      i2<=x"0003";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0003";
      i2<=x"0003";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0003";
      i2<=x"0003";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0001";
      i1<=x"0003";
      i2<=x"0003";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0000";
      i2<=x"0000";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0000";
      i2<=x"0000";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0000";
      i2<=x"0000";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0000";
      i2<=x"0000";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0000";
      i2<=x"0001";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0000";
      i2<=x"0001";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0000";
      i2<=x"0001";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0000";
      i2<=x"0001";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0000";
      i2<=x"0002";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0000";
      i2<=x"0002";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0000";
      i2<=x"0002";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0000";
      i2<=x"0002";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0000";
      i2<=x"0003";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0000";
      i2<=x"0003";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0000";
      i2<=x"0003";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0000";
      i2<=x"0003";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0001";
      i2<=x"0000";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0001";
      i2<=x"0000";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0001";
      i2<=x"0000";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0001";
      i2<=x"0000";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0001";
      i2<=x"0001";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0001";
      i2<=x"0001";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0001";
      i2<=x"0001";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0001";
      i2<=x"0001";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0001";
      i2<=x"0002";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0001";
      i2<=x"0002";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0001";
      i2<=x"0002";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0001";
      i2<=x"0002";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0001";
      i2<=x"0003";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0001";
      i2<=x"0003";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0001";
      i2<=x"0003";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0001";
      i2<=x"0003";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0002";
      i2<=x"0000";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0002";
      i2<=x"0000";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0002";
      i2<=x"0000";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0002";
      i2<=x"0000";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0002";
      i2<=x"0001";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0002";
      i2<=x"0001";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0002";
      i2<=x"0001";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0002";
      i2<=x"0001";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0002";
      i2<=x"0002";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0002";
      i2<=x"0002";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0002";
      i2<=x"0002";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0002";
      i2<=x"0002";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0002";
      i2<=x"0003";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0002";
      i2<=x"0003";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0002";
      i2<=x"0003";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0002";
      i2<=x"0003";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0003";
      i2<=x"0000";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0003";
      i2<=x"0000";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0003";
      i2<=x"0000";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0003";
      i2<=x"0000";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0003";
      i2<=x"0001";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0003";
      i2<=x"0001";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0003";
      i2<=x"0001";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0003";
      i2<=x"0001";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0003";
      i2<=x"0002";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0003";
      i2<=x"0002";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0003";
      i2<=x"0002";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0003";
      i2<=x"0002";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0003";
      i2<=x"0003";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0003";
      i2<=x"0003";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0003";
      i2<=x"0003";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0002";
      i1<=x"0003";
      i2<=x"0003";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0000";
      i2<=x"0000";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0000";
      i2<=x"0000";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0000";
      i2<=x"0000";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0000";
      i2<=x"0000";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0000";
      i2<=x"0001";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0000";
      i2<=x"0001";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0000";
      i2<=x"0001";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0000";
      i2<=x"0001";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0000";
      i2<=x"0002";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0000";
      i2<=x"0002";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0000";
      i2<=x"0002";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0000";
      i2<=x"0002";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0000";
      i2<=x"0003";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0000";
      i2<=x"0003";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0000";
      i2<=x"0003";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0000";
      i2<=x"0003";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0001";
      i2<=x"0000";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0001";
      i2<=x"0000";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0001";
      i2<=x"0000";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0001";
      i2<=x"0000";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0001";
      i2<=x"0001";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0001";
      i2<=x"0001";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0001";
      i2<=x"0001";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0001";
      i2<=x"0001";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0001";
      i2<=x"0002";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0001";
      i2<=x"0002";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0001";
      i2<=x"0002";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0001";
      i2<=x"0002";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0001";
      i2<=x"0003";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0001";
      i2<=x"0003";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0001";
      i2<=x"0003";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0001";
      i2<=x"0003";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0002";
      i2<=x"0000";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0002";
      i2<=x"0000";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0002";
      i2<=x"0000";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0002";
      i2<=x"0000";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0002";
      i2<=x"0001";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0002";
      i2<=x"0001";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0002";
      i2<=x"0001";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0002";
      i2<=x"0001";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0002";
      i2<=x"0002";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0002";
      i2<=x"0002";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0002";
      i2<=x"0002";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0002";
      i2<=x"0002";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0002";
      i2<=x"0003";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0002";
      i2<=x"0003";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0002";
      i2<=x"0003";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0002";
      i2<=x"0003";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0003";
      i2<=x"0000";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0003";
      i2<=x"0000";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0003";
      i2<=x"0000";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0003";
      i2<=x"0000";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0003";
      i2<=x"0001";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0003";
      i2<=x"0001";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0003";
      i2<=x"0001";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0003";
      i2<=x"0001";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0003";
      i2<=x"0002";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0003";
      i2<=x"0002";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0003";
      i2<=x"0002";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0003";
      i2<=x"0002";
      i3<=x"0003";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0003";
      i2<=x"0003";
      i3<=x"0000";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0003";
      i2<=x"0003";
      i3<=x"0001";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0003";
      i2<=x"0003";
      i3<=x"0002";
      wait for 5ns;
      i0<=x"0003";
      i1<=x"0003";
      i2<=x"0003";
      i3<=x"0003";

    end process;
  end;
